Description:    Concept of class inheritance with example 
************************************************************************/
//ADD_CODE: Write a class called parent with property "x" of type int and intialized to 5
//          write a task printf inside the class parent to display the message " THIS IS PARENT CLASS "




//ADD_CODE: Write a class called subclass which is extended from class parent. 
//          Write a task printf inside the class subclass to display the message " THIS IS SUBCLASS "    



    
program inherit;
    
 initial
   begin
//ADD_CODE: Declare handle "p" for class parent and handle "s" for class subclass
    

//ADD_CODE: Create object for handles "p" and "s"
     

//ADD_CODE: Using "s" object access variable "x" and change it's value to 10
     

//ADD_CODE: Display value of "x" using objects "p" and "s" 
     

//ADD_CODE: Call the task printf using objects "p" and "s" 
     

   end
endprogram
